module main

import time

fn (app App) add_activity(user_id int, name string) {
	activity := Activity{
		user_id: user_id
		name: name
		created_at: time.now()
	}

	sql app.db {
		insert activity into Activity
	}
}

fn (mut app App) find_activities(user_id int) []Acti