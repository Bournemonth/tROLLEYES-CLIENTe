module git

pub fn parse_branch_name_from_receive_upload(upload string) ?string {
	uplo