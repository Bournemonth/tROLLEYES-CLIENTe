module main

im