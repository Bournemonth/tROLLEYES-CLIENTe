module main

fn (mut app App) add_star(repo_id