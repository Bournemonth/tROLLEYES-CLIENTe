module main

fn (app App) get_all_repo_branch_nam