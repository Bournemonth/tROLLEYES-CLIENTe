module main

import vweb
import valida