module git

import 