
module main
