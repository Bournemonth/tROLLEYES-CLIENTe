module main

import time

stru