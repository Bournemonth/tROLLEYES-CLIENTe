module main

import ti