
module api

pub struct ApiBranchCount {
	ApiResponse
pub:
	result int
}