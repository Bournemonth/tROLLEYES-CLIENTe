module main

import time

// now only for commits
struct FeedIte