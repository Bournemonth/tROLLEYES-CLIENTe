module highlight

fn init_c() Lang {
	return Lang{
		name: 'C'
		lang_extensions: ['c']
		line_comments: '//'
	