module main

import os

const (
	default_avatar_name  