module main

import rand
import crypto.rand as crypto_rand
import encoding.ba