module config

import os
import json

pub struct Config {
pub:
	repo_storage_path string
	archive_path      string
	avatars_path