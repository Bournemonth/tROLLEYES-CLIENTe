module main

fn (mut app App) watch_repo(repo_id int, user_id int) {
	watch := Watch{
		re