module api

pu