module highlight

fn init_js() Lang {
	return Lang{
		nam